// Class: test_package::test_class
//
// Some description
class test_class;

endclass

// Class: test_package::inherited_class
//
// Some description
class inherited_class extends test_class;

endclass
